`include "pbit.v"
`include "systems.v"

// This module is the top row HA-gates in the sparse multiplier
// Offset of top_row is always assumed to be zero.
module top_row

endmodule

module middle_row

endmodule

module bottom_row

endmodule
